module TopGlove (
    input clk,
    input rst
);
    // TODO
    always @* begin
        
    end
    
endmodule : TopGlove