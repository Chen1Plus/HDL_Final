module TopReceiver (
    input clk,
    input rst
);
    // TODO
endmodule : TopReceiver