module Top (
    input clk,
    input rst
);
    // TODO
endmodule : Top